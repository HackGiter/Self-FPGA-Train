`ifndef __SPM_HEADER__
    `define __SPM_HEADER__
        
    `define SPM_SIZE        16384       //THE CAPACITY OF SPM
    `define SPM_DEPTH       4096        //THE DEPTH OF SPM
    `define SPM_ADDR_W      12          //THE WIDTH OF ADDRESS
    `define SpmAddrBus      11:0        //THE ADDRESS OF BUS
    `define SpmAddrLoc      11:0        //THE LOCATION OF ADDRESS
    
    
`endif 