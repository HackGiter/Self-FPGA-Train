`ifndef __ROM_HEADER__
    `define __ROM_HEADER__
    
    `define ROM_SIZE        8192    //THE SIZE OF ROM
    `define ROM_DEPTH       2048    //THE DEPTH OF ROM
    `define ROM_ADDR_W      11      //THE WIDTH OF ADDRESS
    `define RomAddrBus      10:0    //THE BUS OF ADDRESS
    `define RomAddrLoc      10:0    //THE LOCATION OF ADDRESS
    
    
`endif